module(output y,input a, b);
  assign y = a & b;
endmodule
