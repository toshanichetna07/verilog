module(output y, input a);
  assign y = ~a;
endmodule
